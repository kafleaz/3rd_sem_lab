module and_gate (a, b, c);// module module_name(input, output)
    input a, b;
    output c;
    and and1(c, a, b);
endmodule