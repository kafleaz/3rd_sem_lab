module nor_gate (a, b, c);// module module_name(input, output)
    input a, b;
    output c;
    nor nor1(c, a, b);
endmodule