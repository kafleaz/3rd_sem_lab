module or_gate (a,b,c); //module(keyword) module_name(identifer)(input,output)
input a,b;
output c;
or or1(c,a,b);
endmodule
