module not_gate (a,c); //module(keyword) module_name(identifer)(input,output)
input a;
output c;
not not1(c,a);
endmodule
